module dcachemem(
);